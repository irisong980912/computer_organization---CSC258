// Part 2 skeleton

module part2
	(
		CLOCK_50,						//	On Board 50 MHz
		// Your inputs and outputs here
        KEY,
        SW,
		// The ports below are for the VGA output.  Do not change.
		VGA_CLK,   						//	VGA Clock
		VGA_HS,							//	VGA H_SYNC
		VGA_VS,							//	VGA V_SYNC
		VGA_BLANK_N,						//	VGA BLANK
		VGA_SYNC_N,						//	VGA SYNC
		VGA_R,   						//	VGA Red[9:0]
		VGA_G,	 						//	VGA Green[9:0]
		VGA_B   						//	VGA Blue[9:0]
	);

	input			CLOCK_50;				//	50 MHz
	input   [9:0]   SW;
	input   [3:0]   KEY;

	// Declare your inputs and outputs here
	// Do not change the following outputs
	output			VGA_CLK;   				//	VGA Clock
	output			VGA_HS;					//	VGA H_SYNC
	output			VGA_VS;					//	VGA V_SYNC
	output			VGA_BLANK_N;				//	VGA BLANK
	output			VGA_SYNC_N;				//	VGA SYNC
	output	[9:0]	VGA_R;   				//	VGA Red[9:0]
	output	[9:0]	VGA_G;	 				//	VGA Green[9:0]
	output	[9:0]	VGA_B;   				//	VGA Blue[9:0]
	
	wire resetn;
	assign resetn = KEY[0];
	
	// Create the colour, x, y and writeEn wires that are inputs to the controller.
	wire [2:0] colour;
	wire [7:0] x;
	wire [6:0] y;
	wire writeEn;

	// Create an Instance of a VGA controller - there can be only one!
	// Define the number of colours as well as the initial background
	// image file (.MIF) for the controller.
	vga_adapter VGA(
			.resetn(resetn),
			.clock(CLOCK_50),
			.colour(colour),
			.x(x),
			.y(y),
			.plot(writeEn),
			/* Signals for the DAC to drive the monitor. */
			.VGA_R(VGA_R),
			.VGA_G(VGA_G),
			.VGA_B(VGA_B),
			.VGA_HS(VGA_HS),
			.VGA_VS(VGA_VS),
			.VGA_BLANK(VGA_BLANK_N),
			.VGA_SYNC(VGA_SYNC_N),
			.VGA_CLK(VGA_CLK));
		defparam VGA.RESOLUTION = "160x120";
		defparam VGA.MONOCHROME = "FALSE";
		defparam VGA.BITS_PER_COLOUR_CHANNEL = 1;
		defparam VGA.BACKGROUND_IMAGE = "black.mif";
			
	// Put your code here. Your code should produce signals x,y,colour and writeEn/plot
	// for the VGA controller, in addition to any other functionality your design may require.
    
		combination (CLOCK_50, resetn, KEY[3], KEY[1], SW[6:0], SW[9:7], x, y, colour, writeEn);
	 
	 endmodule
	 
	 
	 //3) combination of datapath and control
	 module combination (CLOCK_50, resetn, go, plot_in, position, colour_in, x, y, colour, writeEn);
		input CLOCK_50, resetn, go, plot_in;
		input [6:0] position;
		input [2:0] colour_in;
		output [7:0] x;
		output [6:0] y;
		output [2:0] colour;
		output plot;
		
		wire ld_x, ld_y, enable;
		
		// control (clk, reset_n, go, plot_in, ld_x, ld_y, plot_out, enable)
		control c0(clk, reset_n, go, plot_in, ld_x, ld_y, plot, enable);
		
		//datapath (clk, enable, reset_n, ld_x, ld_y, position, colour, x_out, y_out, colour_out);
		datapath d0(clk, enable, reset_n, ld_x, ld_y, position, colour, x_out, y_out, colout_out);
	 
	 endmodule
	 
	 
	 
	 
	 
    // Instansiate datapath
	// datapath d0(...);
	module datapath (clk, enable, reset_n, ld_x, ld_y, position, colour, x_out, y_out, colour_out);
		input clk, enable, reset_n, ld_x, ld_y;
		input [6:0] position; // short of switch so only use the first 128 pixels
		input [2:0] colour;
		output [7:0] x_out;
		output [6:0] y_out;
		output [2:0] colour_out;
		
		reg [7:0] x;
		reg [6;0] y;
		reg [2:0] colour;
		
		// loading positions and colour
		always @(posedge clk)
		begin
			if (reset_n == 0)
				begin
					x <= 8'd0;
					y <= 7'd0;
					colour <= 3'd0;
				end
			else
				begin
					x <= ld_x ? {1'b0, position} : x;
					y <= ld_y ? position : y;
					colour <= colour_in;
				end
		end
		
		// counter for a 4x4 square, counting along each row
		reg [3:0] square;
		always @(posedge clk)
		begin
			if (reset_n == 0)
				square <= 4'd0;
			else if (enable)
				begin
					if (square == 4'b1111)
						square <= 4'd0;
					else
						square <= square + 1'b1;
				end
		end
		
		assign x_out = x + square[1:0];
		assign y_out = y + square[3:2];
	
	
	endmodule

	

	
	
    // Instansiate FSM control
    // control c0(...);
	 
	 module control (clk, reset_n, go, plot_in, ld_x, ld_y, plot_out, enable);
			input clk, reset_n, go, plot;
			output ld_x, ld_y, plot_out, enable;
			
			// state table, template given by lab6
			localparam LOAD_X       = 3'd0,
						  LOAD_X_WAIT  = 3'd1,
						  LOAD_Y       = 3'd2,
						  LOAD_Y_WAIT  = 3'd3,
						  PLOT_READY	= 3'd4,
						  PLOT         = 3'd5;
						 
			reg [2:0] current_state, next_state; 
			
			always @(*)
			begin
				case (current_state)
					LOAD_X: next_state = go ? LOAD_X_WAIT : LOAD_X;
					LOAD_X_WAIT: next_state = go ? LOAD_X_WAIT : LOAD_Y;
					LOAD_Y: next_state = go ? LOAD_Y_WAIT : LOAD_Y;
					LOAD_Y_WAIT: next_state = go ? LOAD_Y_WAIT : PLOT_READY;
					PLOT_READY: next_state = plot_in ? PLOT : PLOT_READY;
					PLOT: next_state = go ? LOAD_X : PLOT;
					default: next_state = LOAD_X;
				endcase
			end
			
			always @(*)
			begin:
				  // By default make all our signals 0
				  ld_x = 1'b0;
				  ld_y = 1'b0;
				  ld_c = 1'b0;
				  enable = 1'b0;
				  plot_out = 1'b0;

				  case (current_state)
						LOAD_X: begin
							 ld_x = 1'b1;
						end
						LOAD_Y: begin
							 ld_Y = 1'b1;
						end
						PLOT: begin
							 plot_out = 1'b1;
							 enable = 1'b1;
						end
				  endcase
			end
			
			// current_state registers
		 always@(posedge clk)
		 begin: state_FFs
			  if(reset_n == 0)
					current_state <= LOAD_X;
			  else
					current_state <= next_state;
		 end // state_FFS
		
	 endmodule
	 
